* NGSPICE file created from univ_sr.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

.subckt univ_sr VGND VPWR clk ctrl[0] ctrl[1] d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7]
+ q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] reset
XFILLER_0_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_66_ net11 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_49_ net17 net16 net18 net8 _18_ _17_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_65_ net11 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ net20 _18_ _17_ _23_ _25_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_64_ net11 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_47_ net17 _21_ net9 _24_ VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_63_ net22 _18_ _17_ _34_ _35_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_46_ net1 net2 VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__xnor2_1
Xoutput12 net12 VGND VGND VPWR VPWR q[0] sky130_fd_sc_hd__buf_2
X_62_ net14 _16_ net4 _24_ VGND VGND VPWR VPWR _35_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_45_ net19 _21_ _16_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput13 net13 VGND VGND VPWR VPWR q[1] sky130_fd_sc_hd__clkbuf_4
X_61_ net12 _16_ _21_ VGND VGND VPWR VPWR _34_ sky130_fd_sc_hd__o21a_1
X_44_ net20 _18_ _21_ _22_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput14 net14 VGND VGND VPWR VPWR q[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_60_ net23 _18_ _17_ _31_ _33_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__o32a_1
X_43_ _17_ net10 _19_ net19 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR q[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_42_ net2 VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput16 net16 VGND VGND VPWR VPWR q[4] sky130_fd_sc_hd__buf_2
XFILLER_0_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_41_ net22 _16_ _17_ _20_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR q[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ _18_ net3 _19_ net12 VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput18 net18 VGND VGND VPWR VPWR q[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput19 net19 VGND VGND VPWR VPWR q[7] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 ctrl[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 ctrl[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_79_ clknet_1_1__leaf_clk _15_ _07_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 d[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_78_ clknet_1_0__leaf_clk net21 _06_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 d[1] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_77_ clknet_1_0__leaf_clk _13_ _05_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 d[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_76_ clknet_1_0__leaf_clk _12_ _04_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_59_ net13 _21_ _19_ _32_ VGND VGND VPWR VPWR _33_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 d[3] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_58_ net1 net2 net15 VGND VGND VPWR VPWR _32_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_75_ clknet_1_0__leaf_clk _11_ _03_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_74_ clknet_1_1__leaf_clk _10_ _02_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
Xinput7 d[4] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_57_ net5 _24_ VGND VGND VPWR VPWR _31_ sky130_fd_sc_hd__and2_1
Xinput10 d[7] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_73_ clknet_1_1__leaf_clk net24 _01_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
X_56_ net25 _18_ _17_ _28_ _30_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__o32a_1
Xinput8 d[5] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
Xinput11 reset VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ _18_ _17_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_72_ clknet_1_1__leaf_clk _08_ _00_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
Xinput9 d[6] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ net14 _21_ _19_ _29_ VGND VGND VPWR VPWR _30_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_38_ net1 VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 net18 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
X_71_ net11 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__inv_2
X_54_ _18_ _17_ net16 VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__and3b_1
X_37_ net2 VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__buf_2
Xhold2 _14_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ net11 VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_53_ net6 _24_ VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36_ net1 VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 net13 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ _27_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 net14 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_51_ net16 net15 net17 net7 _18_ _17_ VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 _09_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_50_ _26_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__clkbuf_1
Xhold6 net15 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_69_ net11 VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__inv_2
X_68_ net11 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_67_ net11 VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

