input wire clk,reset,
input wire [1:0]ctrl,
input wire [7:0]d,
output wire [7:0]q);

reg [7:0]r_reg, r_next;

always@(posedge clk, posedge reset)
	if(reset)
	r_reg<=0;
	else
	r_reg<=r_next;

//next_stage logic
always@*
	case(ctrl)
		2'b00: r_next=r_reg; //no operation
		2'b01: r_next={r_reg[6:0], d[0]}; //shift left
		2'b10: r_next={d[7], r_reg[7:1]}; //shift right
		default: r_next=d; //load
	endcase
	
//output logic
assign q=r_reg;
endmodule

		
